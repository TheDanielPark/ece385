version https://git-lfs.github.com/spec/v1
oid sha256:26bb9ec9d654e3e44ec0160eeb6e0c1ed09aa67465368b59a31b7f01f02c5be9
size 542
