module datapath (//input logic Clk, Reset, LD_MDR, LD_MAR, LD_IR, LD_PC, 


);

endmodule

